/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 */
 
package mult_pkg;
typedef enum bit[2:0] {
    RST_OP      	= 3'b000,
    VALID_A_B		= 3'b001,
    INVALID_A_B  	= 3'b010,
    VALID_A_INVALID_B 	= 3'b011,
    VALID_B_INVALID_A 	= 3'b100
} operation_t;

`include "coverage.svh"
`include "tpgen.svh"
`include "scoreboard.svh"
`include "testbench.svh"

endpackage : mult_pkg
