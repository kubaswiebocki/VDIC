/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 */
class maxmult_sequence extends uvm_sequence #(sequence_item);
    `uvm_object_utils(maxmult_sequence)

//------------------------------------------------------------------------------
// local variables
//------------------------------------------------------------------------------

// not necessary, req is inherited
//    sequence_item req;

//------------------------------------------------------------------------------
// constructor
//------------------------------------------------------------------------------

    function new(string name = "maxmult_sequence");
        super.new(name);
    endfunction : new
    
//------------------------------------------------------------------------------
// the sequence body
//------------------------------------------------------------------------------

    task body();
        `uvm_info("SEQ_MAXMULT", "", UVM_MEDIUM)
//      req = sequence_item::type_id::create("req");
//      start_item(req);
//      req.op = mul_op;
//      req.A = 8'hFF;
//      req.B = 8'hFF;
//      finish_item(req);
        `uvm_do_with(req, {op == mul_op; A == 8'hFF; B == 8'hFF;})
        `uvm_do_with(req, {op == rst_op;} )
        `uvm_do_with(req, {op == mul_op;} )
        `uvm_do_with(req, {op == mul_op;} )
        `uvm_do_with(req, {op == rst_op;} )
    endtask : body
    

endclass : maxmult_sequence
